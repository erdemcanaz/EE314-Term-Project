library verilog;
use verilog.vl_types.all;
entity clock_module_vlg_vec_tst is
end clock_module_vlg_vec_tst;
