module fulltemplate (templatey,templatex);

output reg [0:639] templatex;
input [10:0] templatey;

always@(templatey) begin
case(templatey)

0: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
1: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
2: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
3: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
4: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
5: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
6: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
9: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
10: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
11 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
12 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
13 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
14 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
15 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
16 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
17 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
18 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
19 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
20 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
21 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
22 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
23 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
24 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
25 : templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

26: templatex=640'b1111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111;
27: templatex=640'b1111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111;
28: templatex=640'b1111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111;
29: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
30: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
31: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
32: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
33: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
34: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
35: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
36: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
37: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
38: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
39: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
40: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
41: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
42: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
43: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
44: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
45: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
46: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
47: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
48: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
49: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
50: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
51: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
52: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
53: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
54: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
55: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
56: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
57: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111100000000011111111111111111111111100000000111111111111111111111111110000000001111111111111111111111111111100000000000111111111111111111111111000000000001111111111111111111100000001111111111111111111110011111111110011111111111111111111111110011111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
58: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111100111110000111111111111111111111000111100011111111111111111111111110001111000011111111111111111111111111100111111111111111111111111111111111001111111111111111111111111110001111100011111111111111111110011111111110011111111111111111111111110011111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
59: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111100111111100011111111111111111110011111111001111111111111111111111110011111110001111111111111111111111111100111111111111111111111111111111111001111111111111111111111111100011111110001111111111111111110011111111110011111111111111111111111110011111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
60: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110011111111111111111111100111111110011111111111111111100111111111000111111111111111111111110011111111000111111111111111111111111100111111111111111111111111111111111001111111111111111111111111100111111111001111111111111111110011111111110011111111111111111111111110011111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
61: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110011111111111111111111100111111110011111111111111111100111111111111111111111111111111111110011111111100111111111111111111111111100111111111111111111111111111111111001111111111111111111111111001111111111111111111111111111110011111111110011111111111111111111111110011111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
62: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111001111111111111111111100111111100111111111111111111000111111111111111111111111111111111110011111111100111111111111111111111111100111111111111111111111111111111111001111111111111111111111111001111111111111111111111111111110011111111110011111111111111111111111110011111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
63: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111001111111111111111111100000000001111111111111111111000111111111111111111111111111111111110011111111100111111111111111111111111100000000001111111111111111111111111000000000011111111111111111001111111111111111111111111111110000000000000011111111111111111111111110011111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
64: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100111111111111111111100011110000111111111111111111000111111111111111111111111111111111110011111111100111111111111111111111111100000000001111111111111111111111111000000000011111111111111111001111110000001111111111111111110000000000000011111111111111111111111110011111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
65: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100111111111111111111100111111110011111111111111111000111111111111111111111111111111111110011111111100111111111111111111111111100111111111111111111111111111111111001111111111111111111111111001111110000001111111111111111110011111111110011111111111111111111111110011111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
66: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111100111111110011111111111111111100111111111111111111111111111111111110011111111100111111111111111111111111100111111111111111111111111111111111001111111111111111111111111001111111111001111111111111111110011111111110011111111111111111111111110011111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
67: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111110011111111111111111100111111110011111111111111111100111111111000111111111111111111111110011111111000111111111111111111111111100111111111111111111111111111111111001111111111111111111111111100111111111001111111111111111110011111111110011111111111111111111111110011111111111111111111111110111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
68: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111001111111111111111100111111110011111111111111111100011111111001111111111111111111111110011111111001111111111111111111111111100111111111111111111111111111111111001111111111111111111111111100011111111001111111111111111110011111111110011111111111111111111111110011111111111111111111111100011111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
69: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111001111111111111111100111111000011111111111111111110001111110011111111111111111111111110011111100011111111111111111111111111100111111111111111111111111111111111001111111111111111111111111110001111110001111111111111111110011111111110011111111111111111111111110011111111111111111111111110001111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
70: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111111111111111100000000001111111111111111111111100000000111111111111111111111111110000000001111111111111111111111111111100000000000011111111111111111111111001111111111111111111111111111100000000011111111111111111110011111111110011111111111111111111111110011111111111111111111111111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
71: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
72: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
73: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
74: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
75: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
76: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
77: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111000000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
78: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111000000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
79: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111000000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
80: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111000000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
81: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111000000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
82: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111000000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
83: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111000000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
84: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111000000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
85: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111000000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
86: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111000000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
87: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111101111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111000000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
88: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
89: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
90: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
91: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
92: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
93: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
94: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
95: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
96: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
97: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
98: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
99: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111110000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
100: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
101: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
102: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
103: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
104: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
105: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
106: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
107: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
108: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
109: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
110: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
111: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
112: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
113: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
114: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
115: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
116: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
117: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
118: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
119: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
120: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
121: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
122: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
123: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
124: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
125: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000111111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
126: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
127: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
128: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
129: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111110000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
130: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111100000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
131: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
132: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
133: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
134: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
135: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
136: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111101111111111111111110111111111111111111100011111111111111111111111111111111111;
137: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111111110000001111111000111111111111111111111111111001111111111111111110111111111111111111100011111111111111111111111111111111111;
138: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111111000011100011111001111111111111111111111111111001111111111111111110111111111111111111100011111111111111111111111111111111111;
139: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111110001111111001111111111111111111111111111111111001111111111111111110111111111111111111100011111111111111111111111111111111111;
140: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111001111111111111110011111111111111111111111111110011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111100011111111000111111111111111111111111111111111001111111111111111110111111111111111111100011111111111111111111111111111111111;
141: templatex=640'b1111111111111111111111111111111110000100000000000000111111111100111111111111111111111111111111111111111111111001111111111111110011111111111111111111111111100111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111100111111111100111000111100100001111000000111111001111110000000111111111100000001111111100011111111111111111111111111111111111;
142: templatex=640'b1111111111111111111111111111111110000111111100111111111111111111111111111111111111111111111111111111111111111001111111111111110011111111111111111111111111001111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111100111111111111111000111100001111100011110001111001111100111100011111111000111100011111100011111111111111111111111111111111111;
143: templatex=640'b1111111111111111111111111111111110000111111100111111111111111111111111111111111111111111111111111111111111111001111111111111110011111111111111111111111110011111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111100111111111111111000111100111111100111111001111001111001111110001111111001111110011111100011111111111111111111111111111111111;
144: templatex=640'b1111111111111111111111111111111110000111111100111111100100011100111110000001111110110000011111110000011011111001111100000011111111110000001111111111111000111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111100111111111111111000111100111111001111111101111001111001111111001111111001111111111111100011111111111111111111111111111111111;
145: templatex=640'b1111111111111111111111111111111110000111111100111111100001111100111100111100111110001111001111100011100011111001111001111001111111100011100011111111110011111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111100111111111111111000111100111111001111111111111001110000000000001111111100001111111111100011111111111111111111111111111111111;
146: templatex=640'b1111111111111111111111111111111110000111111100111111100111111100111001111110011110011111100111001111110011111001110011111100111111100111110011111111100010000000111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111100111111111111111000111100111111001111111111111001110000000000001111111111000000111111100011111111111111111111111111111111111;
147: templatex=640'b1111111111111111111111111111111110000111111100111111100111111100111111111110011110011111100111001111110011111001110011111100111111100111111111111111100000000000111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111100111111111100111000111100111111001111111111111001110001111111111111111111111100011111100011111111111111111111111111111111111;
148: templatex=640'b1111111111111111111111111111111110000111111100111111100111111100111110000000011110011111100111001111110011111001100000000000111111110000011111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111110011111111000111000111100111111000111111101111001111001111111111111111011111110011111100011111111111111111111111111111111111;
149: templatex=640'b1111111111111111111111111111111110000111111100111111100111111100111000111110011110011111100111001111110011111001100011111111111111111110000111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111111000001111111111111111111111111111111100011111111111110001111110001111000111100111111100111111001111001111000111111011111111001111110011111100011111111111111111111111111111111111;
150: templatex=640'b1111111111111111111111111111111110000111111100111111100111111100111001111110011110011111100111001111110011111001110011111111111111111111110011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000001111111111111111111111111100000011111111111111111111111111111000000111111111111111111111111111111000011111111111111100000000011111000111100111111110000000011111001111100000000011111111100000000111111100011111111111111111111111111111111111;
151: templatex=640'b1111111111111111111111111111111110000111111100111111100111111100111001111100011110011111100111001111110011111001110011111111111111001111110011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111000011111111101111111111111111100001111111101111111100001111111111111000011111111100011111111111111111111111111111111111;
152: templatex=640'b1111111111111111111111111111111110000111111100111111100111111100111000111000011110011111100111100011000011111001111000111000111111100011100011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
153: templatex=640'b1111111111111111111111111111111110000111111100111111100111111100111100000110011110011111100111110000010011111001111100000011111111110000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
154: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
155: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111101111110011111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
156: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
157: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
158: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
159: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
160: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
161: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011110001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
162: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
163: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
164: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
165: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
166: templatex=640'b1111111111111111111111111111111110000100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
167: templatex=640'b1111111111111111111111111111111110000111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
168: templatex=640'b1111111111111111111111111111111110000111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111001111111100111111100111100100001100110000011111111111111111111111100011111111111111111111111111111111111;
169: templatex=640'b1111111111111111111111111111111110000111111100111111101111111011111011001110111000111111111111111111111111111111111111111111111111111111111111111111111111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111001111111100111111100111100000011100000110001111111111111111111111100011111111111111111111111111111111111;
170: templatex=640'b1111111111111111111111111111111110000111111100111111100111111001110000001100000000001111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111001111111100111111100111100011111100011111100111111111111111111111100011111111111111111111111111111111111;
171: templatex=640'b1111111111111111111111111111111110000111111100111111100111111001110001111110011111001111111111111111111111111111111111111111111111111111111111111111100011110001111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111001111111100111111100111100111111100111111100111111111111111111111100011111111111111111111111111111111111;
172: templatex=640'b1111111111111111111111111111111110000111111100111111100111111001110011111110111111101111111111111111111111111111111111111111111111111111111111111111111000000111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111001111111100111111100111100111111100111111100111111111111111111111100011111111111111111111111111111111111;
173: templatex=640'b1111111111111111111111111111111110000111111100111111100111111001110011111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111001111111100111111100111100111111100111111100111111111111111111111100011111111111111111111111111111111111;
174: templatex=640'b1111111111111111111111111111111110000111111100111111100111111001110011111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111001111111100111111100111100111111100111111100111111111111111111111100011111111111111111111111111111111111;
175: templatex=640'b1111111111111111111111111111111110000111111100111111100111111001110011111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111100000001111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111100000001111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111001111111100111111100111100111111100111111100111111111111111111111100011111111111111111111111111111111111;
176: templatex=640'b1111111111111111111111111111111110000111111100111111100111111001110011111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111001111111100011111000111100111111100111111100111111111111111111111100011111111111111111111111111111111111;
177: templatex=640'b1111111111111111111111111111111110000111111100111111100011110001110011111110111111101111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000111111110000000000111100111111100111111100111111111111111111111100011111111111111111111111111111111111;
178: templatex=640'b1111111111111111111111111111111110000111111100111111110000000001110001111100011111000111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111001111111111000001100111100111111100111111100111111111111111111111100011111111111111111111111111111111111;
179: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
180: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
181: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
182: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
183: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
184: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
185: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
186: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
187: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
188: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
189: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111000000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
190: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
191: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011110011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
192: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
193: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111110011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111111000000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
194: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111111100011111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111;
195: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111111100011111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111;
196: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
197: templatex=640'b1111111111111111111111111111111110000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110011111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
198: templatex=640'b1111111111111111111111111111111110000111111111100011111111111111110111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
199: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000111111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
200: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
201: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
202: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
203: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
204: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100001111111111111111111111111111100000001111111111111111111111101010000001000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
205: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111100000001111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
206: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
207: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
208: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
209: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
210: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
211: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110000000000111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
212: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111000000000111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
213: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110011111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
214: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110011111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
215: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110010000111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
216: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110000000001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
217: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111000111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
218: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111100111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
219: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111100111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
220: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110111111100111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
221: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110011111000111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
222: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110001110001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
223: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111100000111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
224: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
225: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
226: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
227: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
228: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
229: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
230: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
231: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111000011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
232: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
233: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000111111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
234: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
235: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
236: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111110000111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
237: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111100011111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
238: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111001111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
239: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110011111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
240: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
241: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100000000011111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
242: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100011111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
243: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111100111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
244: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111100111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
245: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111100111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000011111111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111111111111111111110011111111111111100011111111111111111111111111111111111;
246: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110011111100111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111;
247: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110001111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111;
248: templatex=640'b1111111111111111111111111111111110000111111111100111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111110001111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111;
249: templatex=640'b1111111111111111111111111111111110000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
250: templatex=640'b1111111111111111111111111111111110000111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
251: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
252: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010111110000000111111111111111111111111111000000011111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
253: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
254: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
255: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
256: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111100000001111111111111111111111111100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
257: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
258: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
259: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
260: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
261: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
262: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101000111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
263: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
264: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
265: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
266: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
267: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
268: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
269: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
270: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
271: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
272: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
273: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
274: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
275: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
276: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
277: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
278: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
279: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
280: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
281: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000001111111111111111111111111110000000111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
282: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111110000000111111111111111111111111111100000011000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
283: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
284: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
285: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
286: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
287: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
288: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
289: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
290: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
291: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
292: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
293: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
294: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
295: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
296: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
297: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
298: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001110001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
299: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
300: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
301: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
302: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
303: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111100000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
304: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
305: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
306: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
307: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
308: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
309: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
310: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
311: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
312: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
313: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
314: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110011111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
315: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
316: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
317: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
318: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
319: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
320: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
321: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
322: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
323: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
324: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
325: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
326: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111110000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
327: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111100000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
328: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111000000111111111111111111111111111110000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
329: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100000011111111111111111111111111110000001111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111111000001111111111111111111111111111100000111111111111111111111111111110000111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
330: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111111111111111100000011111111111111111111111111110000000111111111111111111111111110000001111111111111111111111111100000011111111111111111111111111110000011111111111111111111111111110000001111111111111111111111111110000001111111111111111111111111111100000111111111111111111111111111111001111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
331: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
332: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
333: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
334: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
335: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
336: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
337: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
338: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
339: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
340: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
341: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
342: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
343: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
344: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
345: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
346: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
347: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
348: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
349: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
350: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
351: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
352: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
353: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
354: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
355: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
356: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
357: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000100011111111111111111111111111111111111;
358: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000100011111111111111111111111111111111111;
359: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111100111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111001111111111111111111111111111111100100011111111111111111111111111111111111;
360: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111100111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
361: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111100111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
362: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111100111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
363: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
364: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
365: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
366: templatex=640'b1111111111111111111111111111111110000111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
367: templatex=640'b1111111111111111111111111111111110000111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
368: templatex=640'b1111111111111111111111111111111110000111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
369: templatex=640'b1111111111111111111111111111111110000111111110000011111111111111110111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111011111111111111111111111111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
370: templatex=640'b1111111111111111111111111111111110000111111110010001111111110000000000111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111110011111111111111111111111111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111100000000111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111100111101111101111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
371: templatex=640'b1111111111111111111111111111111110000111111100111001111111111111001111111111111111110011111111111111110111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111101111110011111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
372: templatex=640'b1111111111111111111111111111111110000111111100111000111111111111001111111100001111100001111110001111110111111111110001111000111111110000111101111110111110001111111100011111101100111111111111111111111111111111100111111111111111111111111111111100111101111111111111111111111100011111111000111111011111110011111111111111111111111111111100011111111111111111111111111111110011111111111111100111111011111100011111111000111111110001111111110001110000011111111011000111111110000111111110001111111110000011101111110000111111111000111110111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
373: templatex=640'b1111111111111111111111111111111110000111111001111100111111111111001111111001100011110011111001100011110111111110001100000110001111100110011100111110111100110011110011000111001100111111111111111111111111111111100111111111111111111111111111111100111100111100111100110011100001000111100111001110011111110011111111111111111111111111111100011111111111111111111111111111110011111111111111101111111011110001100111100011001111001100011100001000111100111111111000110001111100110011111001100011100111001111101111000110011110000110011110011111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
374: templatex=640'b1111111111111111111111111111111110000111110001111100011111111111001111110111111011110011111111111011110111111110011111001111001111011111101110111100111011111001110111110111111100111111111111111111111111111111100111111111111111111111111111111100111110111000111101110011100111110111101111101111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111100111110011110111110011101111100110011111011100111110111101111111111001111101111011111101110011111011100111101111101111011111001110011111001111111111100111111111111111111111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
375: templatex=640'b1111111111111111111111111111111110000111110011111110011111111111001111100111111001110011111111110011110111111110011111011111101110011111100110011101110011111001110011111111111100111111111111111111111111111111100111111111111111111111111111111100111110111010011001110011100111110111100111111111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111100000001111100111110011001111111110011111011100111110111100111111111001111100110011111100111001111111100111101111101110011111100110011111001111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
376: templatex=640'b1111111111111111111111111111111110000111100011111110001111111111001111100111111001110011111000010011110111111110011111011111001110011111100111011001110000000001111100001111111100111111111111111111111111111111100111111111111111111111111111111100111110011011011011110011100111110111111000011111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111100111001111100000000011001111111110000000011100111110111100111111111001111100110011111100111100000111100111101111101110011111100110011111001111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
377: templatex=640'b1111111111111111111111111111111110000111100111111111001111111111001111100111111001110011110011111011110111111110011111011111101110011111100111001011110011111111111111100111111100111111111111111111111111111111100111111111111111111111111111111100111111010111001011110011100111110111111111001111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111101111100111100111111111001111111110111111111100111110111100111111111001111100110011111100111111110011100111101111101110011111100110011111001111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
378: templatex=640'b1111111111111111111111111111111110000111000111111111100111111111001111110111111011110011110011110011110111111110011111011111101111011111101111100011111011111111110111110011111100111111111111111111111111111111100111111111111111111111111111111100111111000111100011110011100111110111101111100111111111110011111111111111111111111111111100011111111111111111111111111111110011111111111111101111110011100111111111101111100110011111111100111110111100111111111001111101111011111101110011111011100111101111101111011111001110011111001111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
379: templatex=640'b1111111111111111111111111111111110000111001111111111100111111111001111111001100011110001110001000011100111111110011111001111001111100110011111100111111000110001110011000111001100111111111111111111111111111111100111111111111111111111111111111100111111000111100111110011100111110111100111001110011111110011111111111111111111111111111110011111111111111111111111111111100011111111111111100111111011110001100111100011001111001110011100111110011100111111111000110001111100110011111001100011100111100111101111000110011110011111001110011111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
380: templatex=640'b1111111111111111111111111111111110000110011111111111110011111111101111111100001111111001111100011011110111111111111111011111101111110000111111111111111110000111111100011111101100111111111111111111111111111111100111111111111111111111111111111100111111101111110111111011111111110111111000111111011111110011111111111111111111111111111110011111111111111111111111111111110011111111111111101111111111111100001111111000111111110001111111111110111110011111111001000111111110000111111100001111111111110011101111110001111111111111011110111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
381: templatex=640'b1111111111111111111111111111111110000110000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100111111111111111111111000000000000111111111111111111111111111111111111111111111111111111110011111111111111111111111111111100011111111111111111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111000111111111111111111111000000000000100011111111111111111111111111111111111;
382: templatex=640'b1111111111111111111111111111111110000110000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000100011111111111111111111111111111111111;
383: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111011111111100011111111111111111111111111111100111111111111111111111111111111111111111111111111111111110000000000000000000000001111111100011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111000111111111111111111111111111111100100011111111111111111111111111111111111;
384: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
385: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
386: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
387: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
388: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
389: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
390: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
391: templatex=640'b1111111111111111111111111111111110000111110000000000111111110000000000011111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111110011111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111101111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
392: templatex=640'b1111111111111111111111111111111110000111000011111100000111111111001111111111111111110011111111111111110111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111100011111111111111101111110011111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
393: templatex=640'b1111111111111111111111111111111110000100001111111111100011111111001111111110011111100011111110011111110111111111111001111100111111111001111111111111111111001111111100011111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111110011111111000111111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111101111111011111100011111111100111111110011111111110011111000111111111111100111111111001111111110011111111111000111111111111001111111111001111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
394: templatex=640'b1111111111111111111111111111111110000000111111111111110001111111001111111001100111100011111001100011110111111110000100000010001111100010011100111110111100110011110001000111001100111111111111111111111111111111100111111111111111111111111111111100111100111100111100110011100001000111100010001110011111110011111111111111111111111111111110011111111111111111111111111111110011111111111111101111111011110000000111100011001111000100111100000000111000111111111000010001111100010011111001100011100110000111101111100110011110000100011110011111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
395: templatex=640'b1111111111111111111111111111111110000001111111111111111000111111001111110011111011110011110011110011100111111110011111001111001111011111001110111100111011111001110111110111111100111111111111111111111111111111100111111111111111111111111111111100111110111000111101110011100111110111101111101111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111100111110011110111110011101111100110011111011100111110111101111111111001111101111001111001110011111011100111101111101111011111001110011111011111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
396: templatex=640'b1111111111111111111111111111111110000011111111111111111110011111001111100111111001110011111000000011110111111110011111011111101110011111100111011001110000000001111000001111111100111111111111111111111111111111100111111111111111111111111111111100111110011011011011110011100111110111110000011111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111100111001111100000000011001111111110000000011100111110111100111111111001111100110011111100111100001111100111101111101110011111100110011111001111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
397: templatex=640'b1111111111111111111111111111111110000011111111111111111110011111001111100111111001110011111000000011110111111110011111011111101110011111100111011001110000000001111000001111111100111111111111111111111111111111100111111111111111111111111111111100111110011011011011110011100111110111110000011111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111100111001111100000000011001111111110000000011100111110111100111111111001111100110011111100111100001111100111101111101110011111100110011111001111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
398: templatex=640'b1111111111111111111111111111111110000111111111111111111110011111001111100111111001110011110011111011110111111110011111011111101110011111100111001011110011111111111111100111111100111111111111111111111111111111100111111111111111111111111111111100111111010011001011110011100111110111111111001111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111101111100111100111111111001111111110111111111100111110111100111111111001111100110011111100111111110011100111101111101110011111100110011111001111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
399: templatex=640'b1111111111111111111111111111111110000111111111111111111110011111001111110111111011110011110011110011110111111110011111011111101111011111101111100011111011111111110111110011111100111111111111111111111111111111100111111111111111111111111111111100111111000111100011110011100111110111101111100111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111101111110011100111111111001111100110011111111100111110111101111111111001111100111011111101110111111011100111101111101111011111101110011111001111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
400: templatex=640'b1111111111111111111111111111111110000111111111111111111110011111001111110001100011110011110001100011100111111110011111001111001111000110001111100111111000111001110011100111101100111111111111111111111111111111100111111111111111111111111111111100111111000111100111110011100111110111100111001111011111110011111111111111111111111111111110011111111111111111111111111111110011111111111111100111110011110011110111100111001111001110011100111110111100111111111000111001111000110001111001110011100111100111101111001110011110011111001110011111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
401: templatex=640'b1111111111111111111111111111111110000011111111111111111110011111101111111100001111111000111100011011110111111110011111011111101111110000111111110111111110000111111000001111101100111111111111111111111111111111100111111111111111111111111111111100111111101111110111111011101111110111110000011111011111110011111111111111111111111111111110011111111111111111111111111111110011111111111111101111111001111100001111111000011111100000111100111110111110011111111001000011111110000111111100001111101111110011101111110000111111011111011110011111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
402: templatex=640'b1111111111111111111111111111111110000011111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
403: templatex=640'b1111111111111111111111111111111110000001111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
404: templatex=640'b1111111111111111111111111111111110000000111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
405: templatex=640'b1111111111111111111111111111111110000100011111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100111111111111111111111111111111100100011111111111111111111111111111111111;
406: templatex=640'b1111111111111111111111111111111110000110000111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111100011111111111111111111111111111000111111111111111111111111111111111111111111111111111111110011111111111111111111111111111110011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111100011111111111111111111111111111000100011111111111111111111111111111111111;
407: templatex=640'b1111111111111111111111111111111110000111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000100011111111111111111111111111111111111;
408: templatex=640'b1111111111111111111111111111111110000111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
409: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
410: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
411: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
412: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
413: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
414: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
415: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
416: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
417: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
418: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
419: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
420: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
421: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
422: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
423: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
424: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
425: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
426: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
427: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
428: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
429: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
430: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
431: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
432: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
433: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
434: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
435: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
436: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
437: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
438: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
439: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
440: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
441: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
442: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
443: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
444: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
445: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
446: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
447: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
448: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
449: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
450: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
451: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
452: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
453: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
454: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
455: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
456: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
457: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
458: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
459: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
460: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
461: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
462: templatex=640'b1111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111;
463: templatex=640'b1111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111;
464: templatex=640'b1111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111;
465: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111110111111111111111111111111111111111011111111111111111111111111111111011111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111101111111111111111111111111111111101111111111111111111111111111111110111111111111111111111111111111110111111111111111111111111111111110111111111111111111111111111111111011111111111111111111111111111111011111111111111111111111111111111011111111111111111111111111111111001111111111111111111111111111111101111111111111111111111111111111111111111;
466: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
467: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
468: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
469: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
470: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
471: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
472: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
473: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
474: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
475: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
476: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
477: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
478: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
479: templatex=640'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
default: templatex=0;
endcase 

end
endmodule 
