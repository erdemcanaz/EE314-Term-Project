module jkff_chatgpt(
  input wire J,
  input wire K,
  input wire RST,
  input wire CLK,
  output reg Q,
  output reg NQ
);

  always @(posedge CLK or posedge RST) begin
    if (RST)
      Q <= 1'b0;
    else if (J && ~K)
      Q <= 1'b1;
    else if (~J && K)
      Q <= 1'b0;
    else if (J && K)
      Q <= ~Q;
		
	 if (RST)
      NQ <= 1'b1;
    else
      NQ <= ~Q;
  end

	
endmodule
