
module testbench();
	reg D, CLK;
	wire Q;
	
	initial
		begin
		
		
		end
endmodule
