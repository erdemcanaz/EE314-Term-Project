library verilog;
use verilog.vl_types.all;
entity horizontal_and_vertical_counter_vlg_sample_tst is
    port(
        clk_25          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end horizontal_and_vertical_counter_vlg_sample_tst;
