library verilog;
use verilog.vl_types.all;
entity horizontal_and_vertical_counter_vlg_vec_tst is
end horizontal_and_vertical_counter_vlg_vec_tst;
