module fulltemplate (templatey,templatex);

output reg [0:639] templatex;
input [10:0] templatey;

always@(templatey) begin
case(templatey)


0:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
1:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
2:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
3:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
4:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
5:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
6:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
8:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
9:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
10:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
11:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
12:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
13:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
14:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
15:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
16:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
17:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
18:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
19:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
20:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
21:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
22:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
23:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
24:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
25:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
26:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
27:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
28:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
29:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
30:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
31:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
32:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
33:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
34:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
35:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
36:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
37:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
38:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
39:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
40:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
41:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
42:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
43:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
44:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
45:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
46:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
47:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111110000000011111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
48:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111100011111000111111111111111111111111111111111111111111111111111110000000011111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
49:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111001001110010011111111111111111111111111111111111111111111111110000000011111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
50:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111011001110111011111111111111111111111111111111111111111111110000001111111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
51:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010000111101100111001111111111111111111111111111111111111111110000000111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
52:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101011100111101100111001111111111111111111111111111111111111111000000011111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
53:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001011100111101101111101111111111111111111111111111111111111100000001111111111111111111111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
54:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011000000111110001111001111111111111111111111111111111111100000011111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
55:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011000110111110001000001111111111111111111111111111111111000001111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
56:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110100000110111110101111001111111111111111111111111111111110000111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
57:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110011101110111100111111011111111111111111111111111111111100001111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
58:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111101110111001111110011111111111111111111111111111111100011111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
59:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100011101110111011111100011111111111111111111111111111111000111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
60:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110011101110110011111100001111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
61:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110011101110110110111001101111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
62:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110011100000100000001011101111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
63:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000110011100000000001100011100011111111111111111111111111000111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
64:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100100110011100110000001110011100000111111111111111111111110001111111111111111111111111111111111111110111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
65:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110010011001101100110011001001100011111111111111111111100011111111111111111111111111111111111111110011111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
66:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110000010011001101110011100011111001111111111111111111000011111111111111111111111111111111111111110011111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
67:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111100010010011011111111100011111100111111111111111111000111111111111111111111111111111111111111110011111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
68:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011001111000000110011111111100001111100111111111111111110001111111111111111111111111111111111111111111011111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
69:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000011110001100111111111001100111110011111111111111100001111111111111111111111111111111111111111111011111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
70:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111001001111111110001100111110011111111111111100011111111111111111111111111111111111111111111011111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
71:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111100011111100000011111100011111111100011100111111011111111111111000111111111111111111111111111111111111111111111001111111111101111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
72:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111001001111100000011111110011111111000011100111111011111111111111000111111111111111111111111111111111111111111111001111111111001111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
73:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011100000001111110111100111111100011101110011111110011001001111111001111111111110001111111111111111111111111111111111111111111111101111111110011111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
74:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111100000001100111100011111111000111110011111100111000011111111001111111111110001111111111111111111111111111111111111111111111101111111110011111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
75:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111110000000111110001111111110111110011111100111100111111111101111111111100011111111111111111111111111111111111111111111111100111111100111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
76:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111110000111111000111111110011111011111101111100111111111101111111111100011111111111111111111111111111111111111111111111100111111100111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
77:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111110011111100011111111001111001111101111110011111111100111111111000111111111111111111111111111111111111111111111111100111111001111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
78:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111000111110001111111101111100111100111111001111111100111111111000111111111111111111111111111111111111111111111111110111110011111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
79:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000001111111110000000000000000000111100011100111111100111111110111111110001111111111111111111111111111111111111111111111111110011100111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
80:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111100000000000111000111110001110011111100111111110111111110001111111111111111111111111111111111111111111111111110011100111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
81:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111110011011000111000111110111111110111111100011111111111111111111111111111111111111111111111111111010001111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
82:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111011111000011100001110011111110111111100011111111111111111111111111111111111111111111111111111000000111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
83:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111011111101001111000110011111100111111000111111111111111111111111111111111111111111111111111111000000001111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
84:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111101111111011111101110011100010011111100111110000111111111111111111111111111111111111111111111111111111001111000001111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
85:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111001111100111001110010011111100111110001111111111111111111111111111111111111111111111111111111001111110000111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
86:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111000111101111101110010011111001111100011111111111111111111111111111111111111111111111111111111001111111100011111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
87:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111100000001111101111011111111001111100011111111111111111111111111111111111111111111111111111111001111111110001111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
88:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111100011111101111011111110011111000111111111111111111111111111111111111111111111111111111111100111111111000111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
89:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111011111111110011111100111110001111111111111111111111111111111111111111111111111111111111100111111111100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
90:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111111111111110011110001111110001111111111111111111111111111111111111111111111111111111111100111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
91:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000110001111111111111111110111100011111110001111111111111111111111111111111111111111111111111111111111110011111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
92:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100110111111111111100111000111111100011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
93:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001110111111111111111111110001111111100011111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
94:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110011011111111111111100011111000000111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
95:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111001111111111111111100111000000000111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
96:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
97:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
98:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111101111110111110000000011111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
99:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111101111110111110000011111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
100:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111101111110111110011111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
101:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111101111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
102:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
103:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
104:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
105:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101111111111111011111111111111111111111111111111111111111111111111111111111111111110000111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
106:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111011111111111111111111111111111111111111111111111111111111111111111111100000011111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
107:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111011111111111111111111111111111111111111111111111111111111111111111111111100000011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
108:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111101111011111101110100000000000000000000000000001111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
109:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111101111000000000000000000000000000000000000000000000000011111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
110:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011001111111111101111000000000000111111111111111111111111111111000000000000011111111111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
111:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111011111111111101111011111111010111111111111111111111111111111111110000000000000011111111111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
112:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011100011111111111101110011111111000110000110001111111111111111111100100000000000000000001111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
113:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111101110011111111010110011100111001111111111111100110011111111111111100000001111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
114:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000110011111111111101110011111111010110111111111111111111111111001111111111111101111111000000001111111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
115:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011110011111111111101110011111111011111111111111111111101111111111111111111111101111111011110000000111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
116:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111110011111111111101110111111111101111111110111110111101111101111111111111111111111111011111110000000111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
117:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111110011111111111111110111111111101110100111110000111101111111111110100011111111111111111111111110000000111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
118:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111110111111111111111100111111111101110001111111110110101111000111101111110000011111111111111110110111000001111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
119:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111110111111111111111100111111111101111111111111111111111111110000011111111111111111111011111111111111110000011111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
120:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111110111111111111011100111111111101111111111111111111111111111111111111111111111111111011111111111111111100000011111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
121:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111100101111111111111101111111111101111111000000111101111111111111111111111111111111111011011111011111111011100000011111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
122:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111100111111111111111001111111111101110111001000011111111111111111000000111111111111111011111111011111111011111100000111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
123:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111111111111111001111111111101110111111111010111111111111111000001111111111111111111111111011111111011111111000000111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
124:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111111111111111001111111111101110111110000110101111111111101111111111101111111111111101111111111111011111111111000000111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
125:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111100111111111111111011111111111101110111111011001111111111111111000001111111111111111111101111101111111011111111111111000001111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
126:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111100111111111111110011111111111101100111111111111011111111111111111111111111111111111111101111101111111011111111111111111000001111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
127:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111100101111111111110011111111111101101111111111111011111111111111111111111111111111111011111111101111111011111111111111111110000011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
128:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111100101111111111110011111111111101101111111111111111111111111111111111111111111111111011111111101111111011111111111111111111100001110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
129:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111100111111111111110111111111111101101111111111111111111111111110111111101111111111111111110111101111111011111111111111111111111000011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
130:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111100111111111111110111111111111101111111111011111111111111111111011111111111111111110111110111101111111011111111111111111111111110001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
131:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111110111111111111110111111111111101111111111111111111111111111111111111111111111111110111110111101111111011111111111111111111111111100110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
132:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111110111111111111110111111111111101111111111111111111111111111111111011111111111111111111111111101111111011111111111111111111111111110011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
133:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111110111111111111110111111111111101111111111111110111111111111111111111111111111111101111111111101111111011111111111111111111111111111001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
134:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111110111111111111110111111111111101111111111111111111111111111111111111111111111111111111111111101111111011111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
135:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111110111111111111110111111111111111111111111111101111111111111011111111111111111111111111111111101111111011111111111111111111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
136:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111110111111111111110111111111111110111001111111101111111111111101111111111111111111101111111111101111111011111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
137:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111110111011111111110111111111111111111110011111001111111111101111111111111111111111101111111111101111111001111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
138:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111110111011111111110111111111111110111111111111001111111111110111111111111111111111111111111111101111111001111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
139:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001110111011111111110111111111111110111111111111001111111111110111111111111111111111011111111111101111111001111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
140:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000110111111111111110111111111111110011111101111001111111111110111111111111111111111011111111111111111111001111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
141:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111110111111111111110011111100111000111111111110111111111111111111110011111111111111111111001111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
142:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111110111111111111110011111111111110011111111110111111111111111111111011111111111011111111001111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
143:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111110011111111111110011111111101111001111001110111111111111111111111111111111111011111111001111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
144:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011101111111110011111111111110011111111101111000011000101111111011111111111101111111111111011111111001111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
145:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111110011111111111110111111111101111110011111000111111111111111111111111111111111011111111001111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
146:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111110011111111111110011111111101011111111111111110111111111111110011111111111111111111111001111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
147:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111110011111111111110011111111101111111101111111111111101111111100111111111111111111111111011111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
148:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111100000000110011111111111111011111111011111111100111111111111111111011111111111111111111111111111011111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
149:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010000000000000000111111111111011111111111111101100000111111111111011111111111111111111110111111110011111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
150:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111100000000000111111111011111111111110111111111110011111110011111111111111111111110111111110011111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
151:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111000001111111011111111111111111100000011111111111011111111111111111111110111111110011111111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
152:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111000111111011111111111111011111111111101111111111111111111111111111110111111110011111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
153:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111110001111111111111111111111111111111111111111111111111111111111111110111111110011111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
154:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111000000011111111111111111100000111111111111111111111111111111111110111111110011111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
155:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111000000011111111111111111110111111111011111111111111111111111110110111111110011111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
156:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111001110111111111111111111111011111111011111111111111111111111110111111111110011110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
157:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111011111111111111111111001111111111111111111111111100111111011111111111111111111111110111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
158:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111001111111111111111111001110111111111111111011111110111100111111111111111111111111110101111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
159:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111001111111111111111111011110111111111111110001111111111101111111111111111111111111110101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
160:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111001111100000000000011011110111111111111110111111111110111111111111111111111111111111101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
161:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110011111111111111111000111111111111111111111111111111111111111111111111111111111111111101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
162:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011110011111111111111111110011111111111111111111111111111111111111111111111111111111111111101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
163:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111110011111111111111111111001111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
164:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111110011111111111111111111001111110111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
165:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111110011111111111111111111001110110111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
166:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111110011111111111111111111001110110111111111111111111111111111111111111111111111111111111101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
167:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111110011111111111111111111001110111111111111111111111111111111111111111111111111111111111101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
168:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111110011111100111111111111001111111111111111111111111111111111111111111111111111111111111101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
169:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111001111100000011111111001111101111111111111111111111111111111111111111111111111111101111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
170:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111001111111110000001111001111001111111111111111111111111111111111111111111111111111101111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
171:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111001111111111111000010011111111111111111111111111111111111111111111111111111111111101111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
172:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111011111111111111111000011111111111111111111111111111111111111111111111111111111111101111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
173:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111011111111111111111100111111101111111111111111111111111111111111111111111111111111101111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
174:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111111111111011111111111111111110111000101111111111111111111111111111111111111111111111111111101101111011111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
175:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011100011111111111111001111111111111111110000010101111111111111111111111111111111111111111111111111111101101111011111111011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
176:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111110011111111111111001111111111111111110001110101111111111111111111111111111111111111111111111111111101101111011111111010000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
177:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100011111111111111001111111111111111110011000101111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
178:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100111111111111111011111111111111111110010011101111111111111111111111111111111111111111111111111111111111111111111111101111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
179:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100111111111111110011111100001111111110000111101111111111111111111111111111111111111111111111111111110110111111111111101111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
180:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111000111111111111110011111111100001111110001111011111111111111111111111111111111111111111111111111111100111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
181:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111000111111111111110011111111111000011110011111011111111111111111111111111111111111111111111111111111100111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
182:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111001111111111111110011111111111111000110111111011111111111111111111111111111111111111111111111111111100111011111111111110111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
183:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111110001111111111111110011111111111111100000111111011111111111111111111111111111111111111111111111111111111111011101111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
184:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111110001111111111111110011111111111111111001111111011111111111111111111111111111111111111111111111111111111111011111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
185:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111110011111111111111111011111111111111111100100000011111111111111111111111111111111111111111111111111111101111101111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
186:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111110011111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111101110111111111111000000011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
187:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111110011111111111111111111011111111111111110011111100111111111111111111111111111111111111111111111111111111111100111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
188:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111110011111111111111111110000111111111111110011111110111111111111111111111111111111111111111111111111111101111110111111111111111001111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
189:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111100011111111111111111110000001111111111110011111110111111111111111111111111111111111111111111111111111101111110011011111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
190:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111100011111111111111111000110000011111111111011111101111111111111111111111111111111111111111111111111111101111110011111111111001111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
191:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111100011111111111111111001111110000000001111011111101111111111111111111111111111111111111111111111111111111111111001101111111100111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
192:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111000011111111111111100011111111000011111111001111011111111111111111111111111111111111111111111111111111110110111001100011111110111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
193:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111001011111111111110001111111011000011111111001111111111111111111111111111111111111111111111111111111111011111011000110001111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
194:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111011001111111111100011111111011001011111111001111111111111111111111111111111111111111111111111111111111011111101100000110011111000111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
195:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111011001111111111000111111111011011001111111001111111111111111111111111111111111111111111111111111111111000111111101000011001111100001111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
196:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111110011100111111111001111111111011011111111110011111111111111111111111111111111111111111111111111111111111100011111111100011100111100000000111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
197:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111110011100111111111101111111111011011111111000111001111111111111111111111111111111111111111111111111111110110001111110110001110011111111000000001111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
198:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111110111110011111111100111111111011011111110000100001111111111111111111111111111111111111111111111111111111111101111110011001111110111111111100000011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
199:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111100111110011111111110111111110011011111000000001101111111111111111111111111111111111111111111111111111111101111111111011111111111001111111111110000011100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
200:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111100111000011111111110111111110011011100001110111111111111111111111111111111111111111111111111111111111111100111111111111111111111110001111111111100001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
201:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111100110000001111111100111111110110000000111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111110111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
202:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111100100111001111111100111111110110000001111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
203:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111100101111100111111100111111110110011111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
204:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111101001111110011111100111111110110011111111111111111111111111111111111111111111111111111111111111111111011110011111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
205:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111101011111111000111100111111110110011111111111111111011111111111111111111111111111111111111111111111111001110011111110011111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
206:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111101011111111100011100111011111110011111111111111000011111111111111111111111111111111111111111111111111010110011111110011111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
207:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111000011111111111000001111011110110011111111111111001011111111111111111111111111111111111111111111111111010111011111111011111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
208:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111000011101111111110001111011111110011111111111110011011111111111111111111111111111111111111111111111111111011011111111001111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
209:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111000010000111111111101111011111110011111111111110111111111111111111111111111111111111111111111111111111011111001111111101111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
210:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111000011000111111111001111011101110111111111111100111111111111111111111111111111111111111111111111111111111111001111111101111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
211:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111000110000111111111001111011101110111111111111101111111111111111111111111111111111111111111111111111111111111101111111100111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
212:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111000011111111111111001111111101110111111111111001111111111111111111111111111111111111111111111111111111111111101111111100111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
213:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111000011111111111111001111111111110111111111111011111111111111111111111111111111111111111111111111111110111111100111111110111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
214:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111001011111111111111001111011111100111111111110011111111111111111111111111111111111111111111111111111110111111100111111110011111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
215:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111001001111111111111001111011111100111111111110111111011111111111111111111111111111111111111111111111110111111100111111110011111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
216:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101000111111111001101111111111111001111011111100111111111110111111011111111111111111111111111111111111111111111111110111111110111111111011111111111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
217:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001010111111111001100111111111110011111111111100111111111100111111001111111111111111111111111111111111111111111111110111111110011111111001111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
218:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011010111111111001110011111111110011111111111100011111111100111111001111111111111111111111111111111111111111111111111111111110011111111001111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
219:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011010111111111001110001111111110011111111111100001111111101111111111111111111111111111111111111111111111111111111101111111110011111111101111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
220:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110110010111111111001101100111111110011111111111001001111111101111111111111111111111111111111111111111111111111111111101111111111011111111100111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
221:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110010111111111001111110001111110011111111111001101111111101111111110111111111111111111111111111111111111111111111011111111111011111111100111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
222:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110010111111111001111111100000000111110111111001100111111001111111110111111111111111111111111111111111111111111111111111111111001111111110111111111111111111111111111100111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
223:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110010111111111001111111100000000111110111111001100111111011111111110111111111111111111111111111111111111111111111111111111111001111111110011111111101111111111111111100111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
224:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001110110111111111001111111001111000111110111111001110111110011111111110111111111111111111111111111111111111111111110111111111111101111111110011111111100111111111111111100111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
225:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110110011111111001111111011111000111111111111000110111110111111111110011111111111111111111111111111111111111111100111111111111100111111111001111111100111111111111111000111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
226:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011110110011111111001111110011110000111111111111000110111110111111111110011111111111111111111111111111111111111111100111111111111100111111111001111111100111111111011111000111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
227:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110110011111111001111100111110001111111111111000110011100111111111110111101111111111111111111111111111111111111110111111111111100111111111101111111100111111111000111001111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
228:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111110110011111111001111100111100001111111111111000110011100111111111110111101111111111111111111111111111111111111010111111111111110111111111101111111110011111111000111001111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
229:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110110011111111001111001111100001111101111110000011011100111111111110111111111111111111111111111111111111111111010111111111111110111111111100111111110011111111000111001111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
230:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111100110011111111001111011011000001111101111110010011011101111111111110111100111111111111111111111111111111111111010011111111111110011111111100111111110011111111000111001111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
231:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111100110011111111001111011011000101111101111110010011011001111111111110111100111111111111111111111111111111111111010011111111111110011111111110111111110011111111000110011111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
232:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111100110011111111001111001110001101111101111110011011001001111111111110111100111111111111111111111111111111110111110011111111111110011111111110111111111011111111000110011111111101111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
233:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111100111011111111011111101110001101111111111110011001001001111111111100111110111111111111111111111111111111110111110011111111111111011111111110011111111001111111100110011111111001111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
234:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111100111011111111001111101110001001111111111110011001101001111111111100111110111111111111111111111111111111110111110011111111111111011111111110011111111001111111100010011111111001111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
235:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111100111011111111001111100110001001111111111110011001100011111111111100111110111111111111111111111111111111111111111001111111111111001111111111011111111001111111100000011111111011111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
236:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111101111011111111001111100110011001111111111110011001100011111111111101111111111111111111111111111111111111111111111001111111111111001111111111011111111001111111100000111111110011111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
237:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111101111011111111001111100110011001111111111110011001100011111111111101111111111111111111111111111111111111111111111001111111111111001111111111001111111100111111100000111111110011111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
238:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111101111011111111001111110110011001111111111110011001100111111111111001111111111111111111111111111111111111111111111001111111111111001111111111001111111100111111110000111111110011111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
239:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111101111011111111001111110100011001111111111110011101100111111111111001111111111111111111111011111111111101111111111001111111111111001111111111001111111100111111110000111111110111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
240:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111101111011111111101111110100011001111111111110011101100111111111111001111111111111111111111011111111111001111111111001111111111111100111111111001111111100111111110001111111110111111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
241:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111001111011111111100111111100111001111111111110011101100111111111110011111111101111111111111110110111011001111111111001111111111111100111111111100111111110011111110001111111100111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
242:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111001111011111111100111111100111001111101111110011101100111111111110011111111111011011111111011111001011001101111111000111111111111100111111111100111111110011111111001111111100111111110011111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
243:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111001111011111111100111111000111001111101111110011001100111111111110011111111110011111111111011011100011001101111111100111111111111100111111111100111111110011111111001111111101111111100011111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
244:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111001111011111111100111111000111001111101111110011001100111111111100111111111110011101111111111011110011001111111111100111111111111100111111111100111111110011111111001111111101111111000111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
245:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111001111011111111100111111001111001111101111110111001100111111111100111111110001111100111111011011111111001111111111100111111111111110011111111100111111111001111111001111111101111111001111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
246:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111001111011111111110111111001111001111101111110111001100111111111101111111100011111110111111011011111111001111111111100111111111111110011111111110111111111001111111000111111001111110011111111111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
247:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111001111011111111110111110001111001111001111110111001100111111111001111111100011111111111111011100111111001111111111100111111111111110011111111110111111111001111111000111111001111100111111111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
248:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111001111011111111110011110011111001111001111110111001100111111111001111111101111101111000011111100111111001111111111100111111111111110011111111110011111111001111111100111111001111100111111111111111111111111000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
249:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111001111001111111110011110011111001111011110100111001101111111110011111111001111101111001101111101111111001111111111100111111111111110001111111110011111111101111111100111111011111001111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
250:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111001111001111111110011100011111001111011111100111001101111111110111111110001111101111101110111100111111101111111111100111111111111110001111111110011111111100111111100111111011111001111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
251:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111001111001111111110011100011111001111011111100111001101111111100111111110001111111111111110111100111111101111111111110011111111111111001111111110011111111100111111100111111011110011111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
252:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111001111001111111110011100111111001111011111100111001101111111001111111100011111111111111111111100111111101111111111110011111111111111001111111111011111111100111111100111110011100111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
253:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111001111001111111110011000111111001110011111101111001101111111001111111100011111111111111111111100111111101111111111110011111111111111001111111111011111111100111111100011110011100111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111;
254:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111001111001111111110011000111111001110111111101111001101111110011111111000111111111111111111111100111111101111111111110011111111111111001111111111011111111110111111100011110011001111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111;
255:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111001111001111111110011001111111001110111111101111001101111110011111111000111111111111111111111100111111101111111111110011111111111111001111111111001111111110011111100011110011001111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111;
256:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111001111001111111110011001111111001100111101001111001101111110111111111000111111111111111111111100111111100111111111110011111111111111000111111111001111111110011111100011110010011111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111;
257:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111001111111111011001111111001101111101001111011101111100111111110000111111111111111111111110111111100111111111110011111111111111100111111111001111111110011111110011110110111111111111111111111111111000011110001111111111111111111111111111111111111111111111111111111111111111111111111111111111;
258:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111101111111111000001111111011101111111001111011101111001111111100000111111111111111111111110111111100111111111110011111111111111100111111111001111111110011111110011110100111111111111111111111110000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111;
259:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111101111111111000001111111011101111111001111011101110011111111100110111111111111111111111110111111100111111111110011111111111111100111111111001111111111011111110011110001111111111111111111111000000010000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111;
260:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111101111111111100011111111011101111111011110011001110011111111001110111111111111111111111110111111100111111111110011111111111111100111111111101111111111001111110011110001111111111111111111100000111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111;
261:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111100111111111100011111110011101111011011110011001100111111110011110011111111111111111111110111111100111111111110011111111111111100111111111101111111111001111110011110011111111111111111111000111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111;
262:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111100111111111100011111110011101111011011110011011001111111100011110011111111111111111111110111111110111111111111011111111111111110111111111101111111111101111110011110011111111111111111110001111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111;
263:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111100111111111110011111110011101111011011110011011001111111000111110011111111111111111111110011111110111111111111011111111111111110011111111101111111111101111110001110111111111111111111100011111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111;
264:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111101111100111111111110011111110111101111111011110011000011111110001111110011111111111111111111110011111110111111111111011111111111111110011111111101111111111101111110001110111111111111111111000111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111;
265:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111110111111111111001111110111111111111011110111000111111100011111111011111111111111111111110011111110011111111111001111111111111110011111111101111111111100111111001111111111111111111110001111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111;
266:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111110111111111111100111110111111110111011110110001111111100111111111011111111111111111111110011111110011111111111001111111111111110011111111100111111111100111111001111111111111111111100011111111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111;
267:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111100111110011111111111110011100111111110110011100110011111111000111111111001111111111111111111110011111110011111111111001111111111111110011111111100111111111110111111001111111111111111111100111111111111111111111111111100000110000001111111111111111111111111111111111111111111111111111111111111111;
268:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111110111111011111111111111000100111111110110011101110011111110000111111111001111111111111111111110011111110011111111111001111111111111110011111111100111111111110011111001111111111111111111000111111111111111111111111111111000111100000111111111111111111111111111111111111111111111111111111111111111;
269:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111110111111001111111111111100000111111110110011101110111111100000111111111001111111111111111111110011111110011111111111001111111111111110011111111100111111111110011111001111111111111111111001111111111111111111111111111111000111100000011111111111111111111111111111111111111111111111111111111111111;
270:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111110111111001111111111111111100111111110110011001110111111000000011111111101111111111111111111110011111111011111111111001111111111111111011111111100111111111111001111000111111111111111110011111111111111111111111111111100001111110000001111111111111111111111111111111111111111111111111111111111111;
271:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111011111100111111111111111101111111110110000011100111110000000011111111100111111111111111111110011111111011111111111001111111111111111001111111110111111111111001111100111111111111111110011111111111111111111111111111000011111111000000111111111111111111111111111111111111111111111111111111111111;
272:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111011111100111111111111111101111111110110001111101111110000000011111111100111111111111111111110011111111011111111111001111111111111111001111111110111111111111001111100111111111111111100011111111111111111111111111110000111111111000000011111111111111111111111111111111111111111111111111111111111;
273:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111001111110111111111111111101111111111110011111001111000101100001111111110111111111111111111110011111111001111111111101111111111111111001111111110111111111111100111100111111111111111100111111111111111111111111111100011111111111110000001111111111111111111111111111111111111111111111111111111111;
274:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111101111110011111111111111001111111111110011111001111001101100001111111110111111111111111111110011111111001111111111101111111111111111001111111110111111111111100111100111111111111111100111111111111111111111111111000011111111111111000000111111111111111111111111111111111111111111111111111111111;
275:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111100111111001111111111111001111111111110011110011110011101100001111111110011111111111111111110011111111001111111111101111111111111111001111111110111111111111100111100011111111111111001111111111111111111111111110001111111111111111100000011111111111111111111111111111111111111111111111111111111;
276:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111100111111001111111111111001111101111110011100111100011101110001111111110011111111111111111110011111111001111111111101111111111111111001111111110111111111111110111110011111111111111001111111111111111111111111100001111111111111111111000000111111111111111111111111111111111111111111111111111111;
277:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111110111111100111111111111001111101111110111100111100111101110000111111111011111111111111111110011111111101111111111101111111111111111001111111110111111111111110111110011111111111111001111111111111111111111111000011111111111111111111110000011111111111111111111111111111111111111111111111111111;
278:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111110011111110011111111111011111101111110111001111000111101110000111111111011111111111111111110011111111101111111111101111111111111111001111111110011111111111110011110011111111111110001111111111111111111111111000111111111111111111111111100000111111111111111111111111111111111111111111111111111;
279:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111011111111001111111111011111101101110010011110000111101111000111111111001111111111111111110011111111101111111111101111111111111111100111111110011111111111111011110001111111111110011111111111111111111111110001111111111111111111111111110000000111111111111111111111111111111111111111111111111;
280:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111001111111001111111111011111101101110000111100110111001111000011111111001111111111111111110011111111101111111111101111111111111111100111111110011111111111111011111001111111111110011111111111111111111111100011111111111111111111111111111100000001111111111111111111111111111111111111111111111;
281:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111100111111100011111110011111111111100011110000110111101111100011111111100111111111111111111011111111100111111111100111111111111111100111111110011111111111111011111001111111111110011111111111111111111111100011111111111111111111111111111111000000011111111111111111111111111111111111111111111;
282:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111100111111111000011110011111111111100111000000100111101111100011111111100111111111111111111011111111100111111111100111111111111111100111111110011111111111111011111001111111111100011111111111111111111111000111111111111111111111111111111111111000001111111111111111111111111111111111111111111;
283:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111110011111111110000000111111011111100110001100100111001111100011111111100111111111111111111011111111100111111111100111111111111111100111111110011111111111111011111100111111111100011111111111111111111110000111111111111111111111111111111111111100000111111111111111111111111111111111111111111;
284:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111001111111111110000111111011111100000011100101111001111100001111111110011111111111111111011111111110111111111100111111111111111100111111110011111111111111001111100111111111100111111111111111111111110001111111111111111111111111111111111111111000001111111111111111111111111111111111111111;
285:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111100011111111111110111111011111100011111100101111001111100001111111110011111111111111111011111111110111111111100111111111111111100111111110011111111111111001111110011111111100111111111111111111111100011111111111111111111111111111111111111111110000111111111111111111111111111111111111111;
286:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111110000111111111110111111111111100011111100101111001111110001111111110011111111111111111011111111110111111111100111111111111111100111111111011111111111111001111110011111111100111111111111111111111100011111111111111111111111111111111111111111111000111111111111111111111111111111111111111;
287:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111100011111111100111111111111100111111101001111001111110001111111111001111111111111111011111111110011111111100111111111111111100111111111011111111111111001111110011111111100111111111111111111111000111111111111111111111111111111111111111111111000011111111111111111111111111111111111111;
288:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111000011111100111111111111100111111101001111001111110000111111111001111111111111111011111111110011111111100111111111111111100111111111011111111111111001111111001111111100111111111111111111111000111111111111111111111111111111111111111111111000001111111111111111111111111111111111111;
289:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111110000001001111111111111100111111001011111001111110000111111111101111111111111111011111111110011111111110111111111111111100111111111011111111111111101111111001111111000111111111111111111110001111111111111111111111111111111111111111100000000000000111111111111111111111111111111111;
290:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111000001111110111111100111111001011111001111110000111111111101111111111111111011111111111011111111110111111111111111100011111111011111111111111101111111000111111000111111111111111111110001111111111111111111111111111111111111100000000000000000001111111111111111111111111111111;
291:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111101111110111111100111111001011111001111110000111111111100111111111111111011111111111001111111110111111111111111100011111111011111111111111101111111100111111000111111111111111111110001111111111111111111111111111111111110000001111111111100000111111111111111111111111111111;
292:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111101111111111111100111111001011111001111111000011111111110111111111111111001111111111001111111110011111111111111110011111111011111111111111101111111100111111000111111111111111111100011111111111111111111111111111111111100001111111111111110000000111111111111111111111111111;
293:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111101111111111111100111111010011111001111111000011111111110011111111111111001111111111001111111110011111111111111110011111111011111111111111101111111110011111000111111111111111111100011111111111111111111111111111111110000111111111111111111100000011111111111111111111111111;
294:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111101111111111111100111111010011111011111111000011111111110011111111111111001111111111101111111110011111111111111110011111111011111111111111101111111110011111000111111111111111111100111111111111111111111111111111111100001111111111111111111110000000111111111111111111111111;
295:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111111111101111101111111100111111010011111011111111000001111111111011111111111111001111111111100111111110011111111111111110011111111011111111111111101111111110011111000111111111111111111000111111111111111111111111111111111000011111111111111111111111000000011111111111111111111111;
296:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111101111111111111100111111010011111011111111100001111111111001111111111111001111111111100111111110011111111111111110011111111011111111111111101111111111001111000111111111111111111000111111111111111111111111111111100001111111111111111111111111100000000111111111111111111111;
297:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111110001111111111111100111110010011111011111111100001111111111001111111111111101111111111110111111111001111111111111110011111111001111111111111001111111111001111000111111111111111111001111111111111111111111111111111100011111111111111111111111111111000000011111111111111111111;
298:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111110001111111111111000111110010011111011111111100000111111111101111111111111101111111111110111111111001111111111111110011111111001111111111111001111111111001111000111111111111111110001111111111111111111111111111111000111111111111111111111111111111100000001111111111111111111;
299:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000001111111111111000001111111111111000111110010011111011111111110000111111111100111111111111100111111111110011111111001111111111111110011111111001111111111111001111111111001111100111111111111111110001111111111111111111111111111110001111111111111111111111111111111110000001111111111111111111;
300:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111100000101111111111111000111110010011111011111111110000011111111100111111111111100111111111111011111111001111111111111110011111111001111111111111001111111111001111100111111111111111110011111111111111111111111111111100011111111111111111111111111111111111100000011111111111111111;
301:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001100000000000001110101111111111111000111110010011111011111111111000001111111110011111111111110111111111111001111111101111111111111111011111111001111111111111011111111111001111100111111111111111110011111111111111111111111111111000011111111111111111111111111111111111111000011111111111111111;
302:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111100000000011110101111111111111000111110110011111011111111111000000111111110011111111111110011111111111001111111101111111111111111011111111001111111111111011111111111001111100111111111111111100011111111111111111111111111111000111111111111111111111111111111111111111100001111111111111111;
303:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111001111100101111111111111001111110110011111011111111111100000011111111011111111111111011111111111101111111100111111111111111001111111001111111111111011111111111001111100011111111111111100011111111111111111111111111110001111111111111111111111111111111111111111110000111111111111111;
304:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111001111100101111111111111001111110110011111011111111111100000001111111001111111111111001111111111100111111100111111111111111001111111001111111111110011111111111001111100011111111111111100011111111111111111111111111110001111111111111111111111111111111111111111111000011111111111111;
305:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111001111100101111111111111001111110110111111011111111111001000000111111101111111111111001111111111100111111110111111111111111001111111001111111111110011111111110001111110011111111111111100111111111111111111111111111100011111111111111111111111111111111111111111111100001111111111111;
306:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111001111100101111111111111001111110110111111011111111111001100000001111101111111111111101111111111110111111110111111111111111001111111001111111111110011111111110001111110011111111111111100111111111111111111111111111000111111111111111111111111111111111111111111111110001111111111111;
307:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111001111100101111111111111001111110110111111011111111111001111000000111100111111111111100111111111110011111110011111111111111001111111001111111111110011111111110001111110011111111111111100111111111111111111111111111000111111111111100111111111111111111111111111111111000111111111111;
308:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111001111100101111111111111001111110110111111011111111111001111100000111110111111111111110111111111111011111110011111111111111001111111001111111111100011111111110001111110011111111111111100111111111111111111111111110001111111111111000111111111111111111111111111111111000011111111111;
309:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111110001111100101111111111111001111110110111111011111111111001111110000011110011111111111110011111111111001111111011111111111111001111111001111111111100111111111110011111110001111111111111000111111111111111111111111110001111111111110001111111111111111111111111111111111100011111111111;
310:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111110001111101101111111111111001111100110111111011111111111001111110000001110011111111111110011111111111001111111001111111111111001111111001111111111100111111111110011111111001111111111111000111111111111111111111111100011111111111100011111111111111111111111111111111111110001111111111;
311:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111110011111101101111111111111001111100110111111011111111111001111110000000111001111111111111001111111111100111111001111111111111001111111001111111111100111111111110011111111001111111111111101111111111111111111111111100111111111111000111111111111111111111111000000001111111001111111111;
312:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111110011111101101111111111111001111100110111111011111111111001111100011100011001111111111111001111111111100111111101111111111111001111111001111111111100111111111110011111111001111111111111111111111111111111111111111100111111111111001111111111111111111111100000000000011111000111111111;
313:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111110011111101100111111111111001111101110111110011111111111001111100111110000100111111111111101111111111110011111100111111111111101111111001111111111000111111111100011111111000111111111111111111111111111111111111111000111111111110011111111111111111111110000001111100000111100111111111;
314:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111110011111101100111111111111001111101100111110011111111111001111100111111000000111111111111100111111111110011111110111111111111100111111001111111111000111111111100011111111100111111111111111111111111111111111111111001111111111100111111111111111111111000001111111111100001100011111111;
315:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111110011111101100111111111111001111101100111110011111111111001111100111111100000011111111111110111111111111011111110011111111111100111111001111111111000111111111100011111111100111111111111111111111111111111111111110001111111111001111111111111111111110000111111111111110000100011111111;
316:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111110011111101100111111111111001111001100111110011111111111001111100111111111000001111111111110011111111111001111110011111111111100111111001111111111001111111111100011111111100111111111111111111111111111111111111110011111111111001111111111111111111100001111111111111111100000011111111;
317:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111110011111101100111111111111001111001100111110011111111111001111100111111111110000011111111110011111111111101111111001111111111100111111001111111111001111111111100000111111100111111111111111111111111111111111111100011111111110011111111111111111111000111111111111111111110000011111111;
318:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110011111001110111111111111001111001100111110011111111111001111100111111111111100000011111111001111111111100111111001111111111100111111001111111111001111111111100000011111100011111111111111111111111111111111111100011111111100111111111111111111110001111111111111111111111100001111111;
319:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110011111001110111111111111001111001100111110011111111111001111100011111111111111000000011111001111111111110111111100111111111100111111001111111111001111111111000000011111110011111111111111111111111111111111111100111111111001111111111111111111000011111111111111111111111110000111111;
320:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110011111001110111111111111001111001100111110011111111111001111100011111111111111110000000001100111111111110011111100111111111100111111001111111111001111111000000110001111110011111111111111111111111111111111111100111111111001111111111111111111000111111111111111111111111110000001111;
321:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110011111001110111111111111000111001100111110011111111111011111111001111111111111111110000000000011111111111001111110011111111100111111011111111111001100000000011110000111110001111111111111111111111111111111111000111111110011111111111111111100001111111111111111111111111111000000001;
322:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110011111001110011111111111100111001100111110011111111111011111111000111111111111111111111000000000000111111001111110011111111110111111001111111110000000000011111110000011111001111111111111111111111111111111111001111111110011111111111111111100011111111111111111111111111111111000000;
323:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110011111001110011111111111100111001100111110011111111111011111111000001111111111111111111111110000000000000000111111011111111110000000000000000000000000111111111110000001111001111111111111111111111111111111111001111111100111111111111111111000111111111111111111111111111111111110000;
324:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110011111001110011111111111100111001101111110011111111111011111111000000111111111111111111111111111000000000000000000001111100000000000011110000000001111111111111110011000011001111111111111111111111111111111110001111111100111111111111111110001111111111111111111111111111111111111110;
325:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110011111001110011111111111100111001101111110011111111111011111110000000011111111111111111111111111111110000000000000000000000000011111111111001111111111111111111110011100000000111111111111111111111111111111110011111111001111111111111111100001111111111111111111111111111111111111111;
326:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111100011111001110011111111111100111001101111110011111111111011111110000000000111111111111111111111111111111111111000000000011111110011111111111001111111111111111111110011110000000111111111111111111111111111111110011111111001111111111111111100011111111111111111111111111111111111111111;
327:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100011111001110011110111101100111011101111110011111111111011111110000011000011111111111111111111111111111111111111111000111111100011111111111101111111111111111111110011111000000111111111111111111111111111111110011111110011111111111111111000111111111111111111111111111111111111111111;
328:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100011111001110011110111101100111011101111110011111111111011111110000011110000111111111111111111111111111111111111111100110000000011111111111101111111111111111111110011111000000111111111111111111111111111111100011111110011111111111111110001111111111111111111111111111111100000111111;
329:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100111111011111011111111101100011011101111110011111111111011111100000111111000000111111111111111111111111111111111111100100110000011111111111101111111111111111110000111111100000001111111111111111111111111111100111111110011111111111111100001111111111111111111111111111111100000000000;
330:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100111111011111001111111101110011011101111110011111111111011111100000111111110000000011111111111111111111111111111111101100111110000011111111100111111111111111000000111111110000001111111111111111111111111111100111111110011111111111111100011111111111111111111111111111111111100000000;
331:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100111111011111001111111100110011011101111110011111111111011111100000111111111100000000000111111111111111111111111111100100111111100000111111100111111111111110000000111111111000000111111111111111111111111111100111111100111111111111111000111111111111111111111111111111111111111111111;
332:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100111111011111001111111100110011011101111110011111111111011111100000111111111110000000000000000111111111111111111111101100111111111000001111100111111111111000001100111111111100000111111111111111111111111111100111111100111111111111111000111111111111111111111111111111111111111111111;
333:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100111111011111001111111110110011011101111110011111111111011111000001111111111100001111000000000000000001111111111111100100111111111111000011100111111111000000111100011111111110000011111111111111111111111111000111111100111111111111110001111111111111111111111111111111111111111111111;
334:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100111111011111101111111111110011011101111110011111111111011111000001111111111100001111111110000000000000000000000000000100111111111111100000100111111000000011111100011111111111000001111111111111111111111111000111111001111111111111110001111111111111111111111111111111111111111111111;
335:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100111111011111101111111111110011011101111110011111111111011111000001111111111100001111111111111110000000000000000000000100111111111111111000000111000000000011111110011111111111000001111111111111111111111111000111111001111111111111100001111111111111111111111111111111111111111111111;
336:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100111111011111101111111111110010011101111110011111111111011111000001111111111000011111111111111111111100000000000000000100111111111111111100000000000001110011111110011111111111100000111111111111111111111111000111111001111111111111100001111111111111111111111011111111111111111111111;
337:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111000111111011111101111111111110010011001111110011111111111011110000011111111111000011111111111111111111111111111100000000110011111111111111111000000000001110001111110001111111111100000111111111111111111111111000111111011111111111111000100111111111111111111111000011111111111111111111;
338:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111000111111011111101111111111110010011001111110011111111111011110000011111111111000011111111111111111111111111111111111110111001111111111111111111000000011111001111110001111111111100000011111111111111111111111000111110011111111111111000110011111111111111111111110000000000011111111111;
339:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111000111111011111101111111111110010011001111110011111111111011110000011111111110000111111111111111111111111111111111111110011100011111111111111111111100011111001111111001111111111100100011111111111111111111111001111110011111111111111001110011111111111111111111111111001110001111111111;
340:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111000111111011111001111111111110010011001111110011111111111011100000011111111110000111111111111111111111111111111111111111000000000111111111111111111000011111000111111001111111111100110001111111111111111111111001111110011111111111110001111011111111111111111111111111011110000111111111;
341:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111001111111011111001111111111110010011001111110011111111111011100000111111111110000111111111111111111111111111111111111111100000000001111111111111110000011111000111111001111111111100110001111111111111111111111001111110011111111111110001111001111111111111111111111111011111000000111111;
342:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111001111111011111001111111111110000011001111110011111111111011100000111111111100001111111111111111111111111111111111111111111111111000011111111111110000011111100111111000111111111100111000111111111111111111110001111110111111111111110011111001111111111000000111111110011111011000000111;
343:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111001111111011111001111111111110000011001111110011111111111011000000111111111100001111111111111111111111111111111111111111111111111100000111111111100000011111100111111100111111111100111000011111111111111111110001111100111111111111100011111101111111111000000001111110011111001100000000;
344:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111001111111011111001111111111110000011001111110011111111111011000000111111111100001111111111111111111111111111111111111111111111111100000000011111100011001111100011111100111111111100111000011111111111111111110001111100111111111111100011111101111111111111100000111110011111001110000110;
345:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111001111111011111001111111111110000011001111100011111111111011000001111111111000011111111111111111111111111111111111111111111111111100111000000001000111001111100011111100111111111100011110001111111111111111110001111100111111111111100011111100111111111111111000011100111111001110000011;
346:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111001111111011111001111111111110000011001111100011111111111011000001111111111000011111111111111111111111111111111111111111111111111100111111000000000111001111110011111100111111111100011110001111111111111111110001111100111111111111100011111100111111111111111100011100111111001110010001;
347:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111001111111011111001111111111110000011001111100011111111111010000001111111111000011111111111111111111111111111111111111111111111111100011111111000001111000111110001111100011111111100011111000111111111111111110001111100111111111111100011111100111111111111111110000001111111001110011001;
348:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111001111111011111001111111111110010011101111100011111111111010000011111111111000011111111111111111111111111111111111111111111111111100011111111100111111100111110001111110011111111100011111000111111111111111110001111100111111111111100111111100111111111111111111000011111111001110011100;
349:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110001111111011111001111111111110010011101111100011111111111000000011111111110000011111111111111111111111111111111111111111111111111100011111111100111111100111111001111110011111111110011111100011111111111111110001111100111111111111100111111100111111111111111111100011111111001110011110;
350:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110001111111011111001111111111110000011101111100011111111111000000011111111110000111111111111111111111111111111111111111111111111111100011111111100111111100011111001111110001111111110011111100001111111111111110001111100111111111111100111111110011111111111111111110001111111001110011110;
351:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110001111111011111001111111111110000011101111100011111111111000000111111111110000111111111111111111111111111111111111111111111111111100011111111100111111100011111000111110001111111110011111110001111111111111110001111100111111111111100111111110011111111111111111111000111111001110011111;
352:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110001111111011111001111111111110000011101111100011111111111000000111111111110000111111111111111111111111111111111111111111111111111100011111111100111111110011111000111111001111111110011111110000111111111111110001111100111111111111100111111110011111111111111111111000111111101110011111;
353:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110011111111011111001111101111100000011101111100111111111111100000111111111100000111111111111111111111111111111111111111111111111111100011111111100111111110001111100111111001111111110011111111000111111111111110000111100111111111111100111111111001111111111111111111100011111100111001111;
354:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110011111111011111001111101111100100111101111100111111111111000000111111111100000111111111111111111111111111111111111111111111111111100011111111100111111110001111100111111000111111110011111111100111111111111110000111100111111111111100111111111100111111111111111111100011111100111001111;
355:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111110011111111011110011111001111100100111101111100111111111111000000111111111100001111111111111111111111111111111111111111111111111111100011111111100111111111001111100011111000111111110011111111100011111111111110000111100111111111111100111111111110001111111111111111100011111100111001111;
356:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111110011111111011110011111001111100100111100111100111111111111000001111111111100001111111111111111111111111111111111111111111111111111100011111111100111111111001111110011111100111111110001111111100001111111111110000111100111111111111100111111111111000011111111111111100011111100111001111;
357:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111110011111111011110011111011111000100111100111100111111111111000001111111111100001111111111111111111111111111111111111111111111111111100011111111100111111111000111110011111100011111110001111111100000111111111110000111100111111111111100011111111111100001111111111111100111111100111001111;
358:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100011111111011110011111011111001100111100111100111111111111000001111111111000001111111111111111111111111111111111111111111111111111100011111111100111111111100111110001111100011111110001111111100000111111111110000111100111111111111100011111111111111100111111111111100111111100111001111;
359:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100011111111011110011111011111001100111100111100111111111110000001111111111000001111111111111111111111111111111111111111111111111111100011111111100111111111100111111001111110011111110001111111100000011111111110000111100111111111111100011111111111111100011111111111000111111100111001111;
360:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100011111111011110011111011111001100111100111100111111111110000011111111111000001111111111111111111111111111111111111111111111111111100011111111100111111111100111111001111110011111110001111111110000001111111110000111100111111111111100011111111111111110001111111111000111111100111001111;
361:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100011111111011100111110011110001100111100111100111111111110000011111111111000011111111111111111111111111111111111111111111111111111100011111111100111111111110011111000111110001111111001111111110011000111111110000111110011111111111100011111111111111111100111111110001111111100111000111;
362:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111100011111111011100111110111110011100111100111100111111111110000011111111111000011111111111111111111111111111111111111111111111111111100011111111100111111111110011111000111110001111111001111111110011000011111110000111110011111111111100011111111111111111100011111110001111111100111000111;
363:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111100011111111011100111110111110011100111100111100111111111110000111111111110000011111111111111111111111111111111111111111111111111111100011111111100111111111110001111100111111001111111001111111110011100001111110000011110011111111111100011111111111111111110011111100011111111100111000111;
364:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111100111111111011001111110111100011100111110111100111111111100000111111111110000011111111111111111111111111111111111111111111111111111100011111111100111111111110001111100111111000111111001111111110001110000111110000011110011111111111100011111111111111111110001111000111111111100011000111;
365:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111100111111111011001111100111100111100111110111100111111111100000111111111110000111111111111111111111111111111111111111111111111111111100011111111100111111111111001111100011111000111111001111111110001111000011111000011110011111111111110011111111111111111111000000001111111111100011100111;
366:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111000111111111011001111101111100111100111110111100111111111100000111111111110000111111111111111111111111111111111111111111111111111111100011111111100111111111111001111100011111100111111001111111111001111100001111000011110001111111111110011111111111111111111100000011111111111100011100111;
367:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111000111111111011001111101111000111100111110111100111111111100000111111111110000111111111111111111111111111111111111111111111111111111100011111111100111111111111000111110011111100011111001111111111001111110000111000011110001111111111110011111111111111111111111111111111111111100011100111;
368:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111000111111111011001111101111000111100111110111100111111111000001111111111100000111111111111111111111111111111111111111111111111111111100011111111100111111111111000111110011111100011111001111111111001111110000111000011111001111111111110001111111111111111111111111111111111111100011100111;
369:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111000111111111011011111001111001111100111110011100111111111000001111111111100000111111111111111111111111111111111111111111111111111111100011111111100111111111111100111110001111100011111000111111111001111111100001000011111001111111111110001111111111111111111111111111111111111110011100111;
370:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111000111111111010011111011111001111100111110011100111111111000001111111111100000111111111111111111111111111111111111111111111111111111100011111111100111111111111100111110001111100001111000111111111001111111110001000011111001111111111110001111111111111111111111111111111111111110011100111;
371:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111000111111111010011111011111001111100111110011100111111111000001111111111100001111111111111111111111111111111111111111111111111111111100011111111100111111111111100011111001111110001111000111111111001111111110000000001111001111111111111001111111111111111111111111111111111111110011100111;
372:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111000111111111010011110011111001111100111110011100111111111000011111111111100001111111111111111111111111111111111111111111111111111111100011111111100111111111111100011111001111110001111100111111111000111111111000000001111000111111111111001111111111111111111111111111111111111110011100011;
373:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111001111111111010011110111110001111100111110011100111111110000011111111111000001111111111111111111111111111111111111111111111111111111100011111111100111111111111110011111000111110001111100111111111100111111111100000001111000111111111111001111111111111111111111111111111111111110011100011;
374:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111001111111111010011110111110011111100111110011100111111110000011111111111000001111111111111111111111111111111111111111111111111111111100011111111100111111111111110011111100111111000111100111111111100111111111110000001111100111111111111000111111111111111111111111111111111111110011100011;
375:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111001111111111010011110111110011111100111110011100111111110000011111111111000001111111111111111111111111111111111111111111111111111111100011111111100111111111111110001111100111111000111100111111111100111111111111000001111100111111111111000111111111111111111111111111111111111110011100011;
376:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111001111111111010011110110110011111100111110011100111111110000011111111111000001111111111111111111111111111111111111111111111111111111100011111111100111111111111110001111100111111000111100111111111100111111111111000001111100111111111111000111111111111111111111111111111111111110011100011;
377:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111001111111110010011111110110011111100111111011100111111110000111111111111000011111111111111111111111111111111111111111111111111111111100011111111100111111111111111001111100111111000011100111111111100111111111111110000111100011111111111100111111111111111111111111111111111111110011100011;
378:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110001111111110010011111110110011111100111111011100111111100000111111111110000011111111111111111111111111111111111111111111111111111111100011111111100111111111111111001111100011111000011100111111111100111111111111110000111100011111111111100111111111111111111111111111111111111110011100011;
379:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110001111111110010011111110110011111100111111011100111111100000111111111110000011111111111111111111111111111111111111111111111111111111100011111111100111111111111111001111100011111100011100111111111100111111111111110000111100011111111111100111111111111111111111111111111111111110011100011;
380:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110001111111110010011111100110011111100111111011100111111100000111111111110000011111111111111111111111111111111111111111111111111111111100011111111100111111111111111000111110011111100011100111111111100011111111111111000011100011111111111100011111111111111111111111111111111111110011110011;
381:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111110001111111110010011111100110011111100111111011100111111100000111111111110000011111111111111111111111111111111111111111111111111111111100011111111100111111111111111000111110011111100011100011111111100011111111111111000011110011111111111100011111111111111111111111111111111111110011110011;
382:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111110001111111110110011111101110011111100111111011100111111100001111111111110000111111111111111111111111111111111111111111111111111111111100011111111100111111111111111100111110001111110001100011111111110011111111111111100011110011111111111110011111111111111111111111111111111111110011100011;
383:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111110001111111110110011111101100011111100111111011100111111000001111111111110000111111111111111111111111111111111111111111111111111111111100011111111110111111111111111100111110001111110001100011111111110011111111111111100001110001111111111110011111111111111111111111111111111111110011100011;
384:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111110001111111110100011111101100011111100111111011100111111000001111111111100000111111111111111111111111111111111111111111111111111111111100011111111110111111111111111100111110001111110001100011111111110011111111111111110001110001111111111110011111111111111111111111111111111111110011100011;
385:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111110011111111110100011111001100111111100111111001100111111000001111111111100000111111111111111111111111111111111111111111111111111111111100011111111110111111111111111100111111001111110001110011111111110011111111111111111000110001111111111110001111111111111111111111111111111111100011100011;
386:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111110011111111110100011111001100111111100111111001100111111000001111111111100000111111111111111111111111111111111111111111111111111111111100011111111110111111111111111100011111001111110001110011111111110011111111111111111000111001111111111110001111111111111111111111111111111111100111100011;
387:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111110011111111110110011111011100111111100111111001100111111000001111111111100000111111111111111111111111111111111111111111111111111111111100011111111110111111111111111100011111000111111000110011111111110011111111111111111100011001111111111111000111111111111111111111111111111111100111100011;
388:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111110011111111110110011111011100111111100111111001100111111000011111111111100001111111111111111111111111111111111111111111111111111111111100011111111110111111111111111110011111000111111000110011111111110011111111111111111110011000111111111111000111111111111111111111111111111111100111100011;
389:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111110011111111110110011111011100111111100111111001100111110000011111111111000001111111111111111111111111111111111111111111111111111111111100011111111110111111111111111110011111100111111000110011111111110001111111111111111110001000111111111111100011111111111111111111111111111111100111100011;
390:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111110011111111110110010111011100111111100111111001100111110000011111111111000001111111111111111111111111111111111111111111111111111111111100011111111110111111111111111110011111100111111000110011111111110001111111111111111111000000111111111111100011111111111111111111111111111111000111100111;
391:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111110011111111110110110111011100111111100111111001100111110000011111111111000001111111111111111111111111111111111111111111111111111111111100011111111110111111111111111110011111100011111000010011111111111001111111111111111111100000011111111111110001111111111111111111111111111111001111100111;
392:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111100011111111110100110111011100111111100111111001100111110000011111111111000001111111111111111111111111111111111111111111111111111111111100011111111110111111111111111110011111100011111100010011111111111001111111111111111111110000011111111111110001111111111111111111111111111110001111100111;
393:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111100011111111110100111111011100111111100111111101100111100000111111111111000011111111111111111111111111111111111111111111111111111111111100011111111110011111111111111110001111110011111100010001111111111001111111111111111111111000011111111111111000111111111111111111111111111110011111100111;
394:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111100011111111110100111111011100111111100111111101100111100000111111111111000011111111111111111111111111111111111111111111111111111111111100011111111110011111111111111110001111110011111100010001111111111001111111111111111111111000011111111111111000011111111111111111111111111100011111000111;
395:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111100011111111110100111111011100111111100111111101000111100000111111111110000011111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111001111110011111100011001111111111001111111111111111111111110001111111111111100001111111111111111111111111000111111000111;
396:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111100111111111100100111111011100111111100111111101000111100000111111111110000011111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111001111110001111100001001111111111000111111111111111111111110000111111111111110000111111111111111111111110000111111001111;
397:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111100111111111100100110011011100111111100111111101001111100000111111111110000011111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111001111110001111110001001111111111000111111111111111111111111000111111111111111000011111111111111111111100001111111001111;
398:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111100111111111100100110011011100111111100111111101001111000001111111111110000011111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111001111111001111110001001111111111000111111111111111111111111100011111111111111100001111111111111111111000011111110001111;
399:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111100111111111100100110011011101111111100111111101001111000001111111111110000111111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111000111111001111110001001111111111000111111111111111111111111110001111111111111110000011111111111111110000111111110011111;
400:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111100111111111100100110011011101111111100111111101001111000001111111111110000111111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111000111111001111110000001111111111100011111111111111111111111110000111111111111111000000111111111111000001111111110011111;
401:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111100111111111101100110011011101111111100111111100001111000001111111111100000111111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111100111111100111110000001111111111100011111111111111111111111111000011111111111111110000000001110000000111111111100111111;
402:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111000111111111101100110011011101111111100111111100001111000011111111111100000111111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111100111111100111110000001111111111100011111111111111111111111111100001111111111111111100000000000000001111111111000111111;
403:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111000111111111101100110011011101111111100111111100001111000011111111111100000111111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111100111111100111111000001111111111100011111111111111111111111111110000111111111111111111100000000001111111111111000111111;
404:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111000111111111101100110011011001111111100111111100001110000011111111111100000111111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111100111111100111111000001111111111100011111111111111111111111111111000111111111111111111111111111111111111111110001111111;
405:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111000111111111101100110011011001111111100111111100001110000011111111111100000111111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111100011111100111111000001111111111100001111111111111111111111111111100001111111111111111111111111111111111111100011111111;
406:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111000111111111101101111011011001111111100111111100001110000011111111111100001111111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111100011111100011111000001111111111100001111111111111111111111111111110000111111111111111111111111111111111111000011111111;
407:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111000111111111101101111011011001111111100111111100001110000011111111111000001111111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111110011111100011111000001111111111110001111111111111111111111111111111000001111111111111111111111111111111110000111111111;
408:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111000111111111101101111011011001111111100111111100001110000011111111111000001111111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111110011111110011111000001111111111110001111111111111111111111111111111100000111111111111111111111111111111100001111111111;
409:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111000111111111101101111111111001111111001111111110001100000111111111111000001111111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111110011111110011111100001111111111110001111111111111111111111111111111111000000111111111111111111111111111000011111111111;
410:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111000111111111101101111111111001111111001111111110001100000111111111111000001111111111111111111111111111111111111111111111111111111111111100011111111110011111111111111111110011111110001111100001111111111110001111111111111111111111111111111111110000000111111111111111111111100001111111111111;
411:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111000111111111101101111111111001111111001111111110001100000111111111111000001111111111111111111111111111111111111111111111111111111111111110011111111110011111111111111111110011111110001111100001111111111110000111111111111111111111111111111111111110000000011111111111110000000011111111111111;
412:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111000111111111101101111111111001111111001111111110001100000111111111111000001111111111111111111111111111111111111111111111111111111111111110011111111110011111111111111111110001111110001111100001111111111110000111111111111111111111111111111111111111110000000001111000000000001111111111111111;
413:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111001111111111101101111111111001111111001111111110001100000111111111111000011111111111111111111111111111111111111111111111111111111111111110011111111110011111111111111111110001111111001111100001111111111110000111111111111111111111111111111111111111111110000000000000000001111111111111111111;
414:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111001111111111101101111111111011111111001111111110001100001111111111110000011111111111111111111111111111111111111111111111111111111111111110011111111110011111111111111111111001111111001111110001111111111111000111111111111111111111111111111111111111111111111000000000111111111111111111111111;
415:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111001111111111101101111111111011111111001111111110001000001111111111110000011111111111111111111111111111111111111111111111111111111111111110011111111110011111111111111111111001111111000111110001111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111;
416:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111001111111111101101111111111011111111001111111110001000001111111111110000011111111111111111111111111111111111111111111111111111111111111110011111111110011111111111111111111001111111000111110001111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111;
417:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111001111111111101101111111111011111111001111111110001000001111111111110000011111111111111111111111111111111111111111111111111111111111111110011111111111011111111111111111111001111111000111110001111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111;
418:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111001111111111101101111111111011111111001111111110001000001111111111110000011111111111111111111111111111111111111111111111111111111111111110011111111111011111111111111111111001111111000111110001111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111;
419:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111001111111111001101111111110011111111001111111111000000011111111111110000011111111111111111111111111111111111111111111111111111111111111110011111111111011111111111111111111001111111100111110001111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111;
420:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111001111111111001101111111110011111111001111111111000000011111111111110000111111111111111111111111111111111111111111111111111111111111111110011111111111011111111111111111111001111111100111111000111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111;
421:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111110001111111111001101111111110011111111001111111111000000011111111111100000111111111111111111111111111111111111111111111111111111111111111110011111111111011111111111111111111001111111100111111000111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111;
422:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110001111111111001101111111110011111111001111111111000000011111111111100000111111111111111111111111111111111111111111111111111111111111111110011111111111001111111111111111111000111111100011111000111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111;
423:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110001111111111001101111111110011111111001111111111000000011111111111100000111111111111111111111111111111111111111111111111111111111111111110011111111111001111111111111111111100111111100011111000111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111;
424:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110001111111111001101111111110011111111001111111111000000011111111111100000111111111111111111111111111111111111111111111111111111111111111110011111111111001111111111111111111100111111100011111000111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111;
425:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110001111111111011001111110110011111111001111111111000000111111111111100001111111111111111111111111111111111111111111111111111111111111111110001111111111001111111111111111111100111111110011111000011111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111;
426:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110001111111111011001111111110011111111001111111111000000111111111111100001111111111111111111111111111111111111111111111111111111111111111110001111111111001111111111111111111100111111110011111000011111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111;
427:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110001111111111011001111111110011111111001111111111100000111111111111100001111111111111111111111111111111111111111111111111111111111111111110001111111111001111111111111111111100111111110011111100011111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111;
428:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110001111111111011001111111110011111111001111111111100000111111111111000001111111111111111111111111111111111111111111111111111111111111111110001111111111001111111111111111111100111111110011111100011111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111;
429:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110001111111111011001111111110011111111001111111111100001111111111111000001111111111111111111111111111111111111111111111111111111111111111111001111111111001111111111111111111100111111110001111100011111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111;
430:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110001111111110011001111111110011111111001111111111000001111111111111000001111111111111111111111111111111111111111111111111111111111111111111001111111111001111111111111111111100011111111001111100011111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111;
431:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110001111111110011001111111100011111111001111111111000001111111111111000001111111111111111111111111111111111111111111111111111111111111111111001111111111001111111111111111111110011111111001111100011111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111;
432:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111110001111111110011001111101100011111111001111111111000001111111111111000001111111111111111111111111111111111111111111111111111111111111111111001111111111001111111111111111111110011111111001111100011111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111;
433:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111110001111111110011001111111100011111111001111111111000011111111111110000011111111111111111111111111111111111111111111111111111111111111111111001111111111001111111111111111111110011111111001111100001111111111110010011111111111111111111111111111111111111111111111111111111111111111111111111111;
434:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111110001111111110011001111111100011111111001111111111000011111111111110000011111111111111111111111111111111111111111111111111111111111111111111001111111111001111111111111111111110011111111001111100001111111111110010011111111111111111111111111111111111111111111111111111111111111111111111111111;
435:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111110001111111110011001111111100011111111001111111110000011111111111110000011111111111111111111111111111111111111111111111111111111111111111111001111111111001111111111111111111110011111111000111110001111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111;
436:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111110001111111110111001111111100011111111001111111110000011111111111110000011111111111111111111111111111111111111111111111111111111111111111111001111111111001111111111111111111110011111111100111110001111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111;
437:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111110001111111110111001111011100011111111001111111110000011111111111110000011111111111111111111111111111111111111111111111111111111111111111111001111111111001111111111111111111110011111111100111110001111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111;
438:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111110001111111110111001111011100011111111001111111110000011111111111110000011111111111111111111111111111111111111111111111111111111111111111111001111111111001111111111111111111110001111111100111110001111111111110001001111111111111111111111111111111111111111111111111111111111111111111111111111;
439:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111110001111111100111001111011100011111111001111111110000011111111111110000011111111111111111111111111111111111111111111111111111111111111111111000111111111001111111111111111111110001111111100111110001111111111111001001111111111111111111111111111111111111111111111111111111111111111111111111111;
440:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111110001111111100111001111011100011111111001111111100000011111111111110000111111111111111111111111111111111111111111111111111111111111111111111000111111111001111111111111111111110001111111100111110001111111111111001001111111111111111111111111111111111111111111111111111111111111111111111111111;
441:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111110001111111100111001111011100011111110001111111100000111111111111100000111111111111111111111111111111111111111111111111111111111111111111111100111111111101111111111111111111111001111111100011111000111111111111001001111111111111111111111111111111111111111111111111111111111111111111111111111;
442:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111110001111111100111001111011100011111110011111111100000111111111111100000111111111111111111111111111111111111111111111111111111111111111111111100111111111101111111111111111111111001111111110011111000111111111111001001111111111111111111111111111111111111111111111111111111111111111111111111111;
443:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
444:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
445:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
446:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
447:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
448:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
449:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
450:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
451:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
452:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
453:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
454:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
455:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
456:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
457:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
458:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
459:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
460:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
461:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
462:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
463:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
464:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
465:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
466:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
467:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
468:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
469:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
470:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
471:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
472:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
473:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
474:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
475:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
476:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
477:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
478:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
479:templatex=640'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;

default: templatex=0;
endcase 

end
endmodule 
