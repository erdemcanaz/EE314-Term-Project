library verilog;
use verilog.vl_types.all;
entity main_vga_module_vlg_vec_tst is
end main_vga_module_vlg_vec_tst;
