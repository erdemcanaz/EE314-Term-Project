library verilog;
use verilog.vl_types.all;
entity tb_clock_module is
end tb_clock_module;
